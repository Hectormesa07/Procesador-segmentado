
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.NUMERIC_STD.all;


entity INSTRUCTION_MEMORY_MODULE is
    Port ( PC : in  STD_LOGIC_VECTOR (5 downto 0);
           RST : in  STD_LOGIC;
           INSTRUCTION : out  STD_LOGIC_VECTOR (31 downto 0));
end INSTRUCTION_MEMORY_MODULE;

architecture IM of INSTRUCTION_MEMORY_MODULE is

	type ROM_TYPE is array (0 to 63) of std_logic_vector (31 downto 0);

	signal ROM: ROM_TYPE := (	"10100000000100000010000000000100", -- mov 4,%l0
"00000000100000000000000000000000", -- nop
"10100010000100000010000000000101", -- mov 5,%l1
"00000000100000000000000000000000", -- nop
"00000000100000000000000000000000", -- nop
"10100000000000000000000000000000", -- mov comp 
"00000000100000000000000000000000", -- nop
"10100010000000000000000000000000", -- mov comp
"00000000100000000000000000000000", -- nop
"10100100000100000010000000000000", -- mov 0,%l2
"00000000100000000000000000000000", -- nop
"10100100000100000010000000000000", -- mov 0,%l3
"00000000100000000000000000000000", -- nop
"00000000100000000000000000000000", -- nop
"10100100000100000010000000000000", -- mov comp
"00000000100000000000000000000000", -- nop
"10100110000100000010000000000000", -- mov comp
"10000000101001000100000000010011", -- subcc %l1,%l3,%g0
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00110010100000000000000000000101", -- bne 
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00110000100000000000000000001101", -- ba 
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"10100110000001001110000000000001", -- add %l3,1,%l3
"00000000100000000000000000000000",
"10101000000001010000000000010000", -- add %l0,%l4,%l4
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"10100110000100000010000000000000", -- mov comp
"00000000100000000000000000000000",
"10101000000100000010000000000000", -- mov comp
"00110000101111111111111111101100", -- ba 
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
"00000000100000000000000000000000",
									 others => "00000000100000000000000000000000");

begin
process(RST,ROM,PC)
	begin
		if(RST = '1') then
			INSTRUCTION<="00000000000000000000000000000000";
		else
			INSTRUCTION<=ROM(TO_integer(UNSIGNED(PC)));
		end if;
end process;

end IM;